// This packge contains parameter definitions

package top_pkg;

// parameter for mac_unit
    localparam DATA_WIDTH = 8;    
    localparam ACC_DATA_WIDTH = (2*DATA_WIDTH);

    
endpackage