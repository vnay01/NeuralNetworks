`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Vinay Singh
// 
// Create Date: 05/18/2023 09:37:06 PM
// Design Name: mem_controller
// Module Name: mem_controller
//////////////////////////////////////////////////////////////////////////////////


module memory_controller(
                        clk,
                        reset,
                        mem_write,
                        mem_read,
                        fifo_status,
                        memory_address,
                        mem_control_signals
//                        memory_full,
//                        memory_empty
                        );
                        
// Port direction
input clk;
input reset;
input mem_write;
input mem_read;
input [1:0]fifo_status;
//input [19:0] data_in;   // input data from FIFO.
output reg [1:0]mem_control_signals;        // en and wea
output reg [9:0] memory_address;    //memory address generated by controller.
//output reg [19:0] data_out; // represents each element of convoluted matrix.
//output reg memory_full;
//output reg memory_empty;                        


// Internal registers and counters
parameter STATE_SIZE = 3;

parameter IDLE=3'b001,
          READ=3'b010,
          WRITE=3'b100;

reg [STATE_SIZE - 1 : 0 ] current_state, next_state;

//wire [19:0] w_data_in;
//reg [63:0] sampling_register;

reg [9_:0] w_memory_address , w_memory_address_next; 
reg ram_en, write_en;



//assign w_data_in = data_in;
// register update

    always@(posedge clk)
        begin
            if(!reset) 
                begin
                current_state <= IDLE;
                w_memory_address <= {10{1'b0}};
                end
                else
                begin
                current_state <= next_state;
                w_memory_address <= w_memory_address_next;
                end     
        end


// State Change logic
    always@(*)    
        begin
            next_state = current_state;
            w_memory_address_next = w_memory_address;   // preserve current address
            ram_en = 1'b0;
            write_en = 1'b0;

            case(current_state)
                
                IDLE: begin
                        ram_en = 1'b0;
                        write_en = 1'b0;
                        
                        if((mem_write) && (fifo_status == 2'b01)) begin
                         // Ensures that the FIFO buffer is emptied first                                
                            next_state = WRITE;
                            end
             
                      if(mem_read)begin
                        next_state = READ;
                        end                        
                    end
                
                READ: begin
                        ram_en = 1'b1;
                        write_en = 1'b0;
//                        if(!memory_empty)
                        w_memory_address_next = w_memory_address - 1;
                        next_state = IDLE;
                      end
                
                WRITE: begin
                         ram_en = 1'b1;
                         write_en = 1'b1;
//                         if(!memory_full)
                         w_memory_address_next = w_memory_address + 1;
                         next_state = IDLE;
                         end
                
                default:  w_memory_address_next = w_memory_address;
                
                endcase
        end

/// Signals to activate based in state    
always@(*)
begin
    memory_address = w_memory_address;
    mem_control_signals = {ram_en, write_en};
    
end




endmodule
